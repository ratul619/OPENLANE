VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sync_fifo_16x16
  CLASS BLOCK ;
  FOREIGN sync_fifo_16x16 ;
  ORIGIN 0.000 0.000 ;
  SIZE 200.000 BY 200.000 ;
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 97.840 10.640 99.440 187.920 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 187.920 ;
    END
    PORT
      LAYER met4 ;
        RECT 174.640 10.640 176.240 187.920 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 26.730 194.360 28.330 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 179.910 194.360 181.510 ;
    END
  END VPWR
  PIN address_to_read[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 136.040 4.000 136.640 ;
    END
  END address_to_read[0]
  PIN address_to_read[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 37.440 200.000 38.040 ;
    END
  END address_to_read[10]
  PIN address_to_read[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 54.440 4.000 55.040 ;
    END
  END address_to_read[11]
  PIN address_to_read[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 142.840 200.000 143.440 ;
    END
  END address_to_read[12]
  PIN address_to_read[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 159.840 4.000 160.440 ;
    END
  END address_to_read[13]
  PIN address_to_read[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 61.240 200.000 61.840 ;
    END
  END address_to_read[14]
  PIN address_to_read[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 12.970 196.000 13.250 200.000 ;
    END
  END address_to_read[15]
  PIN address_to_read[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 138.550 0.000 138.830 4.000 ;
    END
  END address_to_read[1]
  PIN address_to_read[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 119.040 200.000 119.640 ;
    END
  END address_to_read[2]
  PIN address_to_read[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 112.240 4.000 112.840 ;
    END
  END address_to_read[3]
  PIN address_to_read[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 17.040 200.000 17.640 ;
    END
  END address_to_read[4]
  PIN address_to_read[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 151.430 0.000 151.710 4.000 ;
    END
  END address_to_read[5]
  PIN address_to_read[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 116.010 0.000 116.290 4.000 ;
    END
  END address_to_read[6]
  PIN address_to_read[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 34.040 4.000 34.640 ;
    END
  END address_to_read[7]
  PIN address_to_read[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 193.290 0.000 193.570 4.000 ;
    END
  END address_to_read[8]
  PIN address_to_read[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 27.240 200.000 27.840 ;
    END
  END address_to_read[9]
  PIN address_to_write[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 170.750 0.000 171.030 4.000 ;
    END
  END address_to_write[0]
  PIN address_to_write[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 154.650 196.000 154.930 200.000 ;
    END
  END address_to_write[10]
  PIN address_to_write[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 144.990 196.000 145.270 200.000 ;
    END
  END address_to_write[11]
  PIN address_to_write[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 146.240 4.000 146.840 ;
    END
  END address_to_write[12]
  PIN address_to_write[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 129.240 200.000 129.840 ;
    END
  END address_to_write[13]
  PIN address_to_write[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 153.040 200.000 153.640 ;
    END
  END address_to_write[14]
  PIN address_to_write[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 170.040 4.000 170.640 ;
    END
  END address_to_write[15]
  PIN address_to_write[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 106.350 0.000 106.630 4.000 ;
    END
  END address_to_write[1]
  PIN address_to_write[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 51.610 0.000 51.890 4.000 ;
    END
  END address_to_write[2]
  PIN address_to_write[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 193.840 4.000 194.440 ;
    END
  END address_to_write[3]
  PIN address_to_write[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 10.240 4.000 10.840 ;
    END
  END address_to_write[4]
  PIN address_to_write[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 122.450 196.000 122.730 200.000 ;
    END
  END address_to_write[5]
  PIN address_to_write[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 35.510 196.000 35.790 200.000 ;
    END
  END address_to_write[6]
  PIN address_to_write[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 41.950 0.000 42.230 4.000 ;
    END
  END address_to_write[7]
  PIN address_to_write[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 80.590 196.000 80.870 200.000 ;
    END
  END address_to_write[8]
  PIN address_to_write[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 186.850 196.000 187.130 200.000 ;
    END
  END address_to_write[9]
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 183.630 0.000 183.910 4.000 ;
    END
  END clk
  PIN data_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 99.910 196.000 100.190 200.000 ;
    END
  END data_in[0]
  PIN data_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 196.510 196.000 196.790 200.000 ;
    END
  END data_in[10]
  PIN data_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 161.090 0.000 161.370 4.000 ;
    END
  END data_in[11]
  PIN data_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 90.250 196.000 90.530 200.000 ;
    END
  END data_in[12]
  PIN data_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 20.440 4.000 21.040 ;
    END
  END data_in[13]
  PIN data_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 51.040 200.000 51.640 ;
    END
  END data_in[14]
  PIN data_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 44.240 4.000 44.840 ;
    END
  END data_in[15]
  PIN data_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 74.840 200.000 75.440 ;
    END
  END data_in[1]
  PIN data_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3.310 196.000 3.590 200.000 ;
    END
  END data_in[2]
  PIN data_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 132.110 196.000 132.390 200.000 ;
    END
  END data_in[3]
  PIN data_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 83.810 0.000 84.090 4.000 ;
    END
  END data_in[4]
  PIN data_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.090 0.000 0.370 4.000 ;
    END
  END data_in[5]
  PIN data_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 122.440 4.000 123.040 ;
    END
  END data_in[6]
  PIN data_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 112.790 196.000 113.070 200.000 ;
    END
  END data_in[7]
  PIN data_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 78.240 4.000 78.840 ;
    END
  END data_in[8]
  PIN data_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 187.040 200.000 187.640 ;
    END
  END data_in[9]
  PIN data_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 67.710 196.000 67.990 200.000 ;
    END
  END data_out[0]
  PIN data_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 19.410 0.000 19.690 4.000 ;
    END
  END data_out[10]
  PIN data_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 9.750 0.000 10.030 4.000 ;
    END
  END data_out[11]
  PIN data_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 176.840 200.000 177.440 ;
    END
  END data_out[12]
  PIN data_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 88.440 4.000 89.040 ;
    END
  END data_out[13]
  PIN data_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 74.150 0.000 74.430 4.000 ;
    END
  END data_out[14]
  PIN data_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 163.240 200.000 163.840 ;
    END
  END data_out[15]
  PIN data_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 3.440 200.000 4.040 ;
    END
  END data_out[1]
  PIN data_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 45.170 196.000 45.450 200.000 ;
    END
  END data_out[2]
  PIN data_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 95.240 200.000 95.840 ;
    END
  END data_out[3]
  PIN data_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 32.290 0.000 32.570 4.000 ;
    END
  END data_out[4]
  PIN data_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 64.490 0.000 64.770 4.000 ;
    END
  END data_out[5]
  PIN data_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 102.040 4.000 102.640 ;
    END
  END data_out[6]
  PIN data_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 108.840 200.000 109.440 ;
    END
  END data_out[7]
  PIN data_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 96.690 0.000 96.970 4.000 ;
    END
  END data_out[8]
  PIN data_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 177.190 196.000 177.470 200.000 ;
    END
  END data_out[9]
  PIN empty
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 164.310 196.000 164.590 200.000 ;
    END
  END empty
  PIN full
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 25.850 196.000 26.130 200.000 ;
    END
  END full
  PIN rd_cs
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 58.050 196.000 58.330 200.000 ;
    END
  END rd_cs
  PIN rd_en
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 128.890 0.000 129.170 4.000 ;
    END
  END rd_en
  PIN rst
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 68.040 4.000 68.640 ;
    END
  END rst
  PIN wr_cs
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 180.240 4.000 180.840 ;
    END
  END wr_cs
  PIN wr_en
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 85.040 200.000 85.640 ;
    END
  END wr_en
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 194.120 187.765 ;
      LAYER met1 ;
        RECT 5.520 9.900 194.120 187.920 ;
      LAYER met2 ;
        RECT 6.990 195.720 12.690 196.000 ;
        RECT 13.530 195.720 25.570 196.000 ;
        RECT 26.410 195.720 35.230 196.000 ;
        RECT 36.070 195.720 44.890 196.000 ;
        RECT 45.730 195.720 57.770 196.000 ;
        RECT 58.610 195.720 67.430 196.000 ;
        RECT 68.270 195.720 80.310 196.000 ;
        RECT 81.150 195.720 89.970 196.000 ;
        RECT 90.810 195.720 99.630 196.000 ;
        RECT 100.470 195.720 112.510 196.000 ;
        RECT 113.350 195.720 122.170 196.000 ;
        RECT 123.010 195.720 131.830 196.000 ;
        RECT 132.670 195.720 144.710 196.000 ;
        RECT 145.550 195.720 154.370 196.000 ;
        RECT 155.210 195.720 164.030 196.000 ;
        RECT 164.870 195.720 176.910 196.000 ;
        RECT 177.750 195.720 186.570 196.000 ;
        RECT 187.410 195.720 190.810 196.000 ;
        RECT 6.990 4.280 190.810 195.720 ;
        RECT 6.990 3.555 9.470 4.280 ;
        RECT 10.310 3.555 19.130 4.280 ;
        RECT 19.970 3.555 32.010 4.280 ;
        RECT 32.850 3.555 41.670 4.280 ;
        RECT 42.510 3.555 51.330 4.280 ;
        RECT 52.170 3.555 64.210 4.280 ;
        RECT 65.050 3.555 73.870 4.280 ;
        RECT 74.710 3.555 83.530 4.280 ;
        RECT 84.370 3.555 96.410 4.280 ;
        RECT 97.250 3.555 106.070 4.280 ;
        RECT 106.910 3.555 115.730 4.280 ;
        RECT 116.570 3.555 128.610 4.280 ;
        RECT 129.450 3.555 138.270 4.280 ;
        RECT 139.110 3.555 151.150 4.280 ;
        RECT 151.990 3.555 160.810 4.280 ;
        RECT 161.650 3.555 170.470 4.280 ;
        RECT 171.310 3.555 183.350 4.280 ;
        RECT 184.190 3.555 190.810 4.280 ;
      LAYER met3 ;
        RECT 4.000 186.640 195.600 187.845 ;
        RECT 4.000 181.240 196.000 186.640 ;
        RECT 4.400 179.840 196.000 181.240 ;
        RECT 4.000 177.840 196.000 179.840 ;
        RECT 4.000 176.440 195.600 177.840 ;
        RECT 4.000 171.040 196.000 176.440 ;
        RECT 4.400 169.640 196.000 171.040 ;
        RECT 4.000 164.240 196.000 169.640 ;
        RECT 4.000 162.840 195.600 164.240 ;
        RECT 4.000 160.840 196.000 162.840 ;
        RECT 4.400 159.440 196.000 160.840 ;
        RECT 4.000 154.040 196.000 159.440 ;
        RECT 4.000 152.640 195.600 154.040 ;
        RECT 4.000 147.240 196.000 152.640 ;
        RECT 4.400 145.840 196.000 147.240 ;
        RECT 4.000 143.840 196.000 145.840 ;
        RECT 4.000 142.440 195.600 143.840 ;
        RECT 4.000 137.040 196.000 142.440 ;
        RECT 4.400 135.640 196.000 137.040 ;
        RECT 4.000 130.240 196.000 135.640 ;
        RECT 4.000 128.840 195.600 130.240 ;
        RECT 4.000 123.440 196.000 128.840 ;
        RECT 4.400 122.040 196.000 123.440 ;
        RECT 4.000 120.040 196.000 122.040 ;
        RECT 4.000 118.640 195.600 120.040 ;
        RECT 4.000 113.240 196.000 118.640 ;
        RECT 4.400 111.840 196.000 113.240 ;
        RECT 4.000 109.840 196.000 111.840 ;
        RECT 4.000 108.440 195.600 109.840 ;
        RECT 4.000 103.040 196.000 108.440 ;
        RECT 4.400 101.640 196.000 103.040 ;
        RECT 4.000 96.240 196.000 101.640 ;
        RECT 4.000 94.840 195.600 96.240 ;
        RECT 4.000 89.440 196.000 94.840 ;
        RECT 4.400 88.040 196.000 89.440 ;
        RECT 4.000 86.040 196.000 88.040 ;
        RECT 4.000 84.640 195.600 86.040 ;
        RECT 4.000 79.240 196.000 84.640 ;
        RECT 4.400 77.840 196.000 79.240 ;
        RECT 4.000 75.840 196.000 77.840 ;
        RECT 4.000 74.440 195.600 75.840 ;
        RECT 4.000 69.040 196.000 74.440 ;
        RECT 4.400 67.640 196.000 69.040 ;
        RECT 4.000 62.240 196.000 67.640 ;
        RECT 4.000 60.840 195.600 62.240 ;
        RECT 4.000 55.440 196.000 60.840 ;
        RECT 4.400 54.040 196.000 55.440 ;
        RECT 4.000 52.040 196.000 54.040 ;
        RECT 4.000 50.640 195.600 52.040 ;
        RECT 4.000 45.240 196.000 50.640 ;
        RECT 4.400 43.840 196.000 45.240 ;
        RECT 4.000 38.440 196.000 43.840 ;
        RECT 4.000 37.040 195.600 38.440 ;
        RECT 4.000 35.040 196.000 37.040 ;
        RECT 4.400 33.640 196.000 35.040 ;
        RECT 4.000 28.240 196.000 33.640 ;
        RECT 4.000 26.840 195.600 28.240 ;
        RECT 4.000 21.440 196.000 26.840 ;
        RECT 4.400 20.040 196.000 21.440 ;
        RECT 4.000 18.040 196.000 20.040 ;
        RECT 4.000 16.640 195.600 18.040 ;
        RECT 4.000 11.240 196.000 16.640 ;
        RECT 4.400 9.840 196.000 11.240 ;
        RECT 4.000 4.440 196.000 9.840 ;
        RECT 4.000 3.575 195.600 4.440 ;
  END
END sync_fifo_16x16
END LIBRARY

