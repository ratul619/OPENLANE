VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO RRAM_ANALOG
  CLASS BLOCK ;
  FOREIGN RRAM_ANALOG ;
  ORIGIN 56.250 20.140 ;
  SIZE 1097.410 BY 1335.730 ;
  PIN ENABLE_WL
    PORT
      LAYER met3 ;
        RECT -30.190 1.345 -0.055 3.375 ;
    END
  END ENABLE_WL
  PIN V1_WL
    PORT
      LAYER met3 ;
        RECT -29.900 21.780 0.165 23.810 ;
    END
  END V1_WL
  PIN V2_WL
    PORT
      LAYER met3 ;
        RECT -29.850 25.130 0.135 27.160 ;
    END
  END V2_WL
  PIN V3_WL
    PORT
      LAYER met3 ;
        RECT -29.820 29.300 0.055 31.330 ;
    END
  END V3_WL
  PIN V4_WL
    PORT
      LAYER met3 ;
        RECT -29.990 34.310 0.145 36.530 ;
    END
  END V4_WL
  PIN IN1_WL[0]
    PORT
      LAYER met3 ;
        RECT -29.750 49.520 0.255 52.170 ;
    END
  END IN1_WL[0]
  PIN IN0_WL[0]
    PORT
      LAYER met3 ;
        RECT -29.780 62.560 0.205 65.210 ;
    END
  END IN0_WL[0]
  PIN IN0_WL[1]
    PORT
      LAYER met3 ;
        RECT -29.840 100.970 0.215 103.620 ;
    END
  END IN0_WL[1]
  PIN IN1_WL[1]
    PORT
      LAYER met3 ;
        RECT -29.760 114.050 -27.110 116.750 ;
    END
  END IN1_WL[1]
  PIN IN1_WL[2]
    PORT
      LAYER met3 ;
        RECT -29.760 120.160 0.165 122.810 ;
    END
  END IN1_WL[2]
  PIN IN0_WL[2]
    PORT
      LAYER met3 ;
        RECT -29.860 133.260 0.125 135.910 ;
    END
  END IN0_WL[2]
  PIN IN0_WL[3]
    PORT
      LAYER met3 ;
        RECT -29.910 171.500 0.205 174.150 ;
    END
  END IN0_WL[3]
  PIN IN1_WL[3]
    PORT
      LAYER met3 ;
        RECT -29.840 184.680 0.155 187.330 ;
    END
  END IN1_WL[3]
  PIN IN1_WL[4]
    PORT
      LAYER met3 ;
        RECT -29.960 190.680 0.095 193.330 ;
    END
  END IN1_WL[4]
  PIN IN0_WL[4]
    PORT
      LAYER met3 ;
        RECT -29.740 203.590 0.245 206.240 ;
    END
  END IN0_WL[4]
  PIN IN0_WL[5]
    PORT
      LAYER met3 ;
        RECT -29.930 242.100 0.045 244.750 ;
    END
  END IN0_WL[5]
  PIN IN1_WL[5]
    PORT
      LAYER met3 ;
        RECT -29.740 255.100 -27.090 257.800 ;
    END
  END IN1_WL[5]
  PIN IN1_WL[6]
    PORT
      LAYER met3 ;
        RECT -29.910 261.210 0.135 263.860 ;
    END
  END IN1_WL[6]
  PIN IN0_WL[6]
    PORT
      LAYER met3 ;
        RECT -29.840 274.390 0.095 277.040 ;
    END
  END IN0_WL[6]
  PIN IN0_WL[7]
    PORT
      LAYER met3 ;
        RECT -29.880 312.770 -27.230 315.470 ;
    END
  END IN0_WL[7]
  PIN IN1_WL[7]
    PORT
      LAYER met3 ;
        RECT -29.930 325.730 0.135 328.380 ;
    END
  END IN1_WL[7]
  PIN IN1_WL[8]
    PORT
      LAYER met3 ;
        RECT -29.840 331.810 0.175 334.460 ;
    END
  END IN1_WL[8]
  PIN IN0_WL[8]
    PORT
      LAYER met3 ;
        RECT -29.790 345.070 0.245 347.720 ;
    END
  END IN0_WL[8]
  PIN IN0_WL[9]
    PORT
      LAYER met3 ;
        RECT -29.960 383.420 0.175 386.070 ;
    END
  END IN0_WL[9]
  PIN IN1_WL[9]
    PORT
      LAYER met3 ;
        RECT -29.840 396.430 0.135 399.080 ;
    END
  END IN1_WL[9]
  PIN IN1_WL[10]
    PORT
      LAYER met3 ;
        RECT -29.810 402.660 0.175 405.310 ;
    END
  END IN1_WL[10]
  PIN IN0_WL[10]
    PORT
      LAYER met3 ;
        RECT -29.860 415.540 0.095 418.190 ;
    END
  END IN0_WL[10]
  PIN IN0_WL[11]
    PORT
      LAYER met3 ;
        RECT -29.880 454.020 0.215 456.670 ;
    END
  END IN0_WL[11]
  PIN IN1_WL[11]
    PORT
      LAYER met3 ;
        RECT -29.960 467.050 -0.035 469.700 ;
    END
  END IN1_WL[11]
  PIN IN1_WL[12]
    PORT
      LAYER met3 ;
        RECT -30.160 473.140 0.045 475.790 ;
    END
  END IN1_WL[12]
  PIN IN0_WL[12]
    PORT
      LAYER met3 ;
        RECT -29.910 486.190 0.175 488.840 ;
    END
  END IN0_WL[12]
  PIN IN0_WL[13]
    PORT
      LAYER met3 ;
        RECT -29.930 524.650 -27.280 527.350 ;
    END
  END IN0_WL[13]
  PIN IN1_WL[13]
    PORT
      LAYER met3 ;
        RECT -30.080 537.600 0.095 540.250 ;
    END
  END IN1_WL[13]
  PIN IN1_WL[14]
    PORT
      LAYER met3 ;
        RECT -29.930 543.790 0.175 546.440 ;
    END
  END IN1_WL[14]
  PIN IN0_WL[14]
    PORT
      LAYER met3 ;
        RECT -30.010 556.870 0.045 559.520 ;
    END
  END IN0_WL[14]
  PIN IN0_WL[15]
    PORT
      LAYER met3 ;
        RECT -29.980 595.270 0.095 597.920 ;
    END
  END IN0_WL[15]
  PIN IN1_WL[15]
    PORT
      LAYER met3 ;
        RECT -29.840 608.480 0.135 611.130 ;
    END
  END IN1_WL[15]
  PIN ENABLE_SL
    PORT
      LAYER met2 ;
        RECT 417.640 -19.210 419.710 210.790 ;
    END
  END ENABLE_SL
  PIN V1_SL
    PORT
      LAYER met2 ;
        RECT 438.060 -19.210 440.330 211.010 ;
    END
  END V1_SL
  PIN V2_SL
    PORT
      LAYER met2 ;
        RECT 441.490 -19.290 443.760 210.980 ;
    END
  END V2_SL
  PIN V3_SL
    PORT
      LAYER met2 ;
        RECT 445.510 -19.290 447.810 -16.850 ;
    END
  END V3_SL
  PIN V4_SL
    PORT
      LAYER met2 ;
        RECT 450.730 -19.210 453.000 210.990 ;
    END
  END V4_SL
  PIN IN1_SL[0]
    PORT
      LAYER met3 ;
        RECT 465.930 -18.880 468.700 211.100 ;
    END
  END IN1_SL[0]
  PIN IN0_SL[0]
    PORT
      LAYER met3 ;
        RECT 478.970 -18.800 481.740 211.050 ;
    END
  END IN0_SL[0]
  PIN IN0_SL[1]
    PORT
      LAYER met3 ;
        RECT 517.190 -19.130 519.960 211.060 ;
    END
  END IN0_SL[1]
  PIN IN1_SL[2]
    PORT
      LAYER met3 ;
        RECT 536.570 -18.960 539.340 211.010 ;
    END
  END IN1_SL[2]
  PIN IN0_SL[2]
    PORT
      LAYER met3 ;
        RECT 549.660 -19.130 552.430 210.970 ;
    END
  END IN0_SL[2]
  PIN IN0_SL[3]
    PORT
      LAYER met3 ;
        RECT 587.800 -18.920 590.570 211.050 ;
    END
  END IN0_SL[3]
  PIN IN1_SL[3]
    PORT
      LAYER met3 ;
        RECT 600.960 -19.040 603.730 211.000 ;
    END
  END IN1_SL[3]
  PIN IN1_SL[4]
    PORT
      LAYER met3 ;
        RECT 606.760 -19.130 609.530 210.940 ;
    END
  END IN1_SL[4]
  PIN IN0_SL[4]
    PORT
      LAYER met3 ;
        RECT 620.140 -18.920 622.910 211.090 ;
    END
  END IN0_SL[4]
  PIN IN0_SL[5]
    PORT
      LAYER met3 ;
        RECT 658.360 -19.040 661.130 210.890 ;
    END
  END IN0_SL[5]
  PIN IN1_SL[5]
    PORT
      LAYER met3 ;
        RECT 671.360 -19.210 674.130 211.080 ;
    END
  END IN1_SL[5]
  PIN IN1_SL[6]
    PORT
      LAYER met3 ;
        RECT 677.610 -19.170 680.380 169.945 ;
    END
  END IN1_SL[6]
  PIN IN0_SL[6]
    PORT
      LAYER met3 ;
        RECT 690.700 -19.040 693.470 210.940 ;
    END
  END IN0_SL[6]
  PIN IN0_SL[7]
    PORT
      LAYER met3 ;
        RECT 728.960 -19.040 731.730 210.980 ;
    END
  END IN0_SL[7]
  PIN IN1_SL[7]
    PORT
      LAYER met3 ;
        RECT 741.800 -19.000 744.570 210.980 ;
    END
  END IN1_SL[7]
  PIN IN1_SL[8]
    PORT
      LAYER met3 ;
        RECT 748.100 -18.880 750.870 211.020 ;
    END
  END IN1_SL[8]
  PIN IN0_SL[8]
    PORT
      LAYER met3 ;
        RECT 761.260 -19.040 764.030 211.090 ;
    END
  END IN0_SL[8]
  PIN IN0_SL[9]
    PORT
      LAYER met3 ;
        RECT 799.780 -19.090 802.550 211.020 ;
    END
  END IN0_SL[9]
  PIN IN1_SL[9]
    PORT
      LAYER met3 ;
        RECT 812.820 -19.290 815.590 210.980 ;
    END
  END IN1_SL[9]
  PIN IN1_SL[10]
    PORT
      LAYER met3 ;
        RECT 818.820 -19.330 821.590 211.020 ;
    END
  END IN1_SL[10]
  PIN IN0_SL[10]
    PORT
      LAYER met3 ;
        RECT 831.950 -18.760 834.720 210.940 ;
    END
  END IN0_SL[10]
  PIN IN0_SL[11]
    PORT
      LAYER met3 ;
        RECT 870.380 -19.210 873.150 211.060 ;
    END
  END IN0_SL[11]
  PIN IN1_SL[11]
    PORT
      LAYER met3 ;
        RECT 883.380 -19.420 886.150 210.810 ;
    END
  END IN1_SL[11]
  PIN IN1_SL[12]
    PORT
      LAYER met3 ;
        RECT 889.470 -19.170 892.240 210.890 ;
    END
  END IN1_SL[12]
  PIN IN0_SL[12]
    PORT
      LAYER met3 ;
        RECT 902.560 -19.170 905.330 211.020 ;
    END
  END IN0_SL[12]
  PIN IN0_SL[13]
    PORT
      LAYER met3 ;
        RECT 940.940 -19.250 943.710 210.890 ;
    END
  END IN0_SL[13]
  PIN IN1_SL[13]
    PORT
      LAYER met3 ;
        RECT 954.105 -18.975 956.715 210.940 ;
    END
  END IN1_SL[13]
  PIN IN0_SL[14]
    PORT
      LAYER met3 ;
        RECT 973.120 -19.000 975.890 210.890 ;
    END
  END IN0_SL[14]
  PIN IN0_SL[15]
    PORT
      LAYER met3 ;
        RECT 1011.670 -19.130 1014.440 210.940 ;
    END
  END IN0_SL[15]
  PIN IN1_SL[15]
    PORT
      LAYER met3 ;
        RECT 1024.800 -19.090 1027.570 210.980 ;
    END
  END IN1_SL[15]
  PIN ENABLE_BL
    PORT
      LAYER met3 ;
        RECT -10.510 927.445 -8.480 1315.590 ;
    END
  END ENABLE_BL
  PIN V1_BL
    PORT
      LAYER met3 ;
        RECT 10.070 927.225 11.870 1315.190 ;
    END
  END V1_BL
  PIN V2_BL
    PORT
      LAYER met3 ;
        RECT 13.425 927.255 15.490 1315.055 ;
    END
  END V2_BL
  PIN V3_BL
    PORT
      LAYER met3 ;
        RECT 17.535 927.335 19.600 1315.305 ;
    END
  END V3_BL
  PIN V4_BL
    PORT
      LAYER met3 ;
        RECT 22.625 927.245 24.690 1315.185 ;
    END
  END V4_BL
  PIN IN1_BL[0]
    PORT
      LAYER met3 ;
        RECT 37.700 927.135 40.300 1315.230 ;
    END
  END IN1_BL[0]
  PIN IN0_BL[0]
    PORT
      LAYER met3 ;
        RECT 50.770 927.185 53.370 1315.300 ;
    END
  END IN0_BL[0]
  PIN IN0_BL[1]
    PORT
      LAYER met3 ;
        RECT 89.100 927.175 91.700 1315.320 ;
    END
  END IN0_BL[1]
  PIN IN1_BL[1]
    PORT
      LAYER met3 ;
        RECT 102.260 927.195 104.860 1315.160 ;
    END
  END IN1_BL[1]
  PIN IN1_BL[2]
    PORT
      LAYER met3 ;
        RECT 108.340 927.225 110.940 1315.200 ;
    END
  END IN1_BL[2]
  PIN IN0_BL[2]
    PORT
      LAYER met3 ;
        RECT 121.420 927.265 124.020 1315.230 ;
    END
  END IN0_BL[2]
  PIN IN0_BL[3]
    PORT
      LAYER met3 ;
        RECT 159.690 927.185 162.290 1315.230 ;
    END
  END IN0_BL[3]
  PIN IN1_BL[3]
    PORT
      LAYER met3 ;
        RECT 172.780 927.235 175.380 1315.060 ;
    END
  END IN1_BL[3]
  PIN IN1_BL[4]
    PORT
      LAYER met3 ;
        RECT 178.890 927.295 181.490 1315.230 ;
    END
  END IN1_BL[4]
  PIN IN0_BL[4]
    PORT
      LAYER met3 ;
        RECT 191.970 927.145 194.570 1315.250 ;
    END
  END IN0_BL[4]
  PIN IN0_BL[5]
    PORT
      LAYER met3 ;
        RECT 230.280 927.345 232.880 1315.330 ;
    END
  END IN0_BL[5]
  PIN IN1_BL[5]
    PORT
      LAYER met3 ;
        RECT 243.430 927.155 246.030 1315.090 ;
    END
  END IN1_BL[5]
  PIN IN1_BL[6]
    PORT
      LAYER met3 ;
        RECT 249.480 927.255 252.080 1315.290 ;
    END
  END IN1_BL[6]
  PIN IN0_BL[6]
    PORT
      LAYER met3 ;
        RECT 262.530 927.295 265.130 1315.220 ;
    END
  END IN0_BL[6]
  PIN IN0_BL[7]
    PORT
      LAYER met3 ;
        RECT 300.830 927.255 303.430 1315.320 ;
    END
  END IN0_BL[7]
  PIN IN1_BL[7]
    PORT
      LAYER met3 ;
        RECT 313.850 927.255 316.450 1315.260 ;
    END
  END IN1_BL[7]
  PIN IN1_BL[8]
    PORT
      LAYER met3 ;
        RECT 320.030 927.215 322.630 1315.190 ;
    END
  END IN1_BL[8]
  PIN IN0_BL[8]
    PORT
      LAYER met3 ;
        RECT 333.190 927.145 335.790 1315.120 ;
    END
  END IN0_BL[8]
  PIN IN0_BL[9]
    PORT
      LAYER met3 ;
        RECT 371.630 927.215 374.230 1315.260 ;
    END
  END IN0_BL[9]
  PIN IN1_BL[9]
    PORT
      LAYER met3 ;
        RECT 384.770 927.255 387.370 1315.230 ;
    END
  END IN1_BL[9]
  PIN IN1_BL[10]
    PORT
      LAYER met3 ;
        RECT 390.830 927.215 393.430 1315.250 ;
    END
  END IN1_BL[10]
  PIN IN0_BL[10]
    PORT
      LAYER met3 ;
        RECT 403.900 927.295 406.500 1315.230 ;
    END
  END IN0_BL[10]
  PIN IN0_BL[11]
    PORT
      LAYER met3 ;
        RECT 442.250 927.175 444.850 1315.250 ;
    END
  END IN0_BL[11]
  PIN IN1_BL[11]
    PORT
      LAYER met3 ;
        RECT 455.370 927.425 457.970 1315.530 ;
    END
  END IN1_BL[11]
  PIN IN1_BL[12]
    PORT
      LAYER met3 ;
        RECT 461.290 927.345 463.890 1315.390 ;
    END
  END IN1_BL[12]
  PIN IN0_BL[12]
    PORT
      LAYER met3 ;
        RECT 474.370 927.215 476.970 1315.250 ;
    END
  END IN0_BL[12]
  PIN IN0_BL[13]
    PORT
      LAYER met3 ;
        RECT 512.870 927.345 515.470 1315.360 ;
    END
  END IN0_BL[13]
  PIN IN1_BL[13]
    PORT
      LAYER met3 ;
        RECT 525.670 927.295 528.270 1315.320 ;
    END
  END IN1_BL[13]
  PIN IN1_BL[14]
    PORT
      LAYER met3 ;
        RECT 531.960 927.215 534.560 1315.300 ;
    END
  END IN1_BL[14]
  PIN IN0_BL[14]
    PORT
      LAYER met3 ;
        RECT 544.990 927.345 547.590 1315.400 ;
    END
  END IN0_BL[14]
  PIN IN0_BL[15]
    PORT
      LAYER met3 ;
        RECT 583.390 927.295 585.990 1315.300 ;
    END
  END IN0_BL[15]
  PIN IN1_BL[15]
    PORT
      LAYER met3 ;
        RECT 596.560 1312.390 599.470 1315.250 ;
    END
  END IN1_BL[15]
  PIN IN1_SL[14]
    PORT
      LAYER met3 ;
        RECT 960.070 -18.960 962.840 211.020 ;
    END
  END IN1_SL[14]
  PIN IN1_SL[1]
    PORT
      LAYER met3 ;
        RECT 530.320 -18.880 533.090 211.040 ;
    END
  END IN1_SL[1]
  PIN CSA[0]
    PORT
      LAYER met2 ;
        RECT 750.995 517.535 1036.590 518.315 ;
    END
  END CSA[0]
  PIN ENABLE_CSA
    PORT
      LAYER met3 ;
        RECT 783.055 725.440 1036.650 729.140 ;
    END
  END ENABLE_CSA
  PIN V0_REF_ADC
    PORT
      LAYER met2 ;
        RECT 817.800 1307.770 819.370 1311.735 ;
    END
  END V0_REF_ADC
  PIN V1_REF_ADC
    PORT
      LAYER met2 ;
        RECT 811.130 1300.500 812.800 1311.375 ;
    END
  END V1_REF_ADC
  PIN V2_REF_ADC
    PORT
      LAYER met2 ;
        RECT 802.130 1291.740 803.640 1311.475 ;
    END
  END V2_REF_ADC
  PIN CSA[1]
    PORT
      LAYER met2 ;
        RECT 750.995 530.575 1036.305 531.465 ;
    END
  END CSA[1]
  PIN CSA[2]
    PORT
      LAYER met2 ;
        RECT 750.995 543.795 1036.105 544.685 ;
    END
  END CSA[2]
  PIN CSA[3]
    PORT
      LAYER met2 ;
        RECT 750.995 556.945 1036.405 557.835 ;
    END
  END CSA[3]
  PIN CSA[4]
    PORT
      LAYER met2 ;
        RECT 750.995 570.055 1036.215 570.945 ;
    END
  END CSA[4]
  PIN CSA[5]
    PORT
      LAYER met2 ;
        RECT 750.995 583.265 1035.625 584.155 ;
    END
  END CSA[5]
  PIN CSA[6]
    PORT
      LAYER met2 ;
        RECT 750.995 596.435 1036.505 597.325 ;
    END
  END CSA[6]
  PIN CSA[7]
    PORT
      LAYER met2 ;
        RECT 750.995 609.525 1036.305 610.415 ;
    END
  END CSA[7]
  PIN CSA[8]
    PORT
      LAYER met2 ;
        RECT 750.995 622.735 1035.505 623.625 ;
    END
  END CSA[8]
  PIN CSA[9]
    PORT
      LAYER met2 ;
        RECT 750.995 635.815 1035.925 636.705 ;
    END
  END CSA[9]
  PIN CSA[10]
    PORT
      LAYER met2 ;
        RECT 750.995 649.095 1034.965 649.985 ;
    END
  END CSA[10]
  PIN CSA[11]
    PORT
      LAYER met2 ;
        RECT 750.995 662.165 1035.835 663.055 ;
    END
  END CSA[11]
  PIN CSA[12]
    PORT
      LAYER met2 ;
        RECT 750.995 675.395 1036.035 676.285 ;
    END
  END CSA[12]
  PIN CSA[13]
    PORT
      LAYER met2 ;
        RECT 750.995 688.505 1036.615 689.395 ;
    END
  END CSA[13]
  PIN CSA[14]
    PORT
      LAYER met2 ;
        RECT 750.995 701.735 1037.135 702.625 ;
    END
  END CSA[14]
  PIN CSA[15]
    PORT
      LAYER met2 ;
        RECT 750.995 714.755 1036.165 715.645 ;
    END
  END CSA[15]
  PIN ADC_OUT0[0]
    PORT
      LAYER met2 ;
        RECT 921.170 741.240 1036.225 742.050 ;
    END
  END ADC_OUT0[0]
  PIN ADC_OUT1[0]
    PORT
      LAYER met2 ;
        RECT 921.115 758.340 1036.035 759.070 ;
    END
  END ADC_OUT1[0]
  PIN ADC_OUT2[0]
    PORT
      LAYER met2 ;
        RECT 919.830 776.850 1035.990 777.610 ;
    END
  END ADC_OUT2[0]
  PIN ADC_OUT0[1]
    PORT
      LAYER met2 ;
        RECT 919.435 802.020 1036.205 802.770 ;
    END
  END ADC_OUT0[1]
  PIN ADC_OUT1[1]
    PORT
      LAYER met2 ;
        RECT 921.010 819.030 1036.060 819.890 ;
    END
  END ADC_OUT1[1]
  PIN ADC_OUT2[1]
    PORT
      LAYER met2 ;
        RECT 921.030 837.610 1036.520 838.470 ;
    END
  END ADC_OUT2[1]
  PIN ADC_OUT0[2]
    PORT
      LAYER met2 ;
        RECT 919.790 862.750 1036.180 863.610 ;
    END
  END ADC_OUT0[2]
  PIN ADC_OUT1[2]
    PORT
      LAYER met2 ;
        RECT 920.060 879.760 1036.510 880.600 ;
    END
  END ADC_OUT1[2]
  PIN ADC_OUT2[2]
    PORT
      LAYER met2 ;
        RECT 919.845 898.360 1036.575 899.170 ;
    END
  END ADC_OUT2[2]
  PIN ADC_OUT0[3]
    PORT
      LAYER met2 ;
        RECT 920.930 923.500 1035.770 924.380 ;
    END
  END ADC_OUT0[3]
  PIN ADC_OUT1[3]
    PORT
      LAYER met2 ;
        RECT 920.410 940.570 1036.300 941.470 ;
    END
  END ADC_OUT1[3]
  PIN ADC_OUT2[3]
    PORT
      LAYER met2 ;
        RECT 919.440 959.170 1036.230 960.030 ;
    END
  END ADC_OUT2[3]
  PIN ADC_OUT0[4]
    PORT
      LAYER met2 ;
        RECT 921.025 984.310 1036.255 985.120 ;
    END
  END ADC_OUT0[4]
  PIN ADC_OUT1[4]
    PORT
      LAYER met2 ;
        RECT 921.130 1001.340 1036.735 1002.150 ;
    END
  END ADC_OUT1[4]
  PIN ADC_OUT2[4]
    PORT
      LAYER met2 ;
        RECT 919.970 1019.930 1036.730 1020.730 ;
    END
  END ADC_OUT2[4]
  PIN ADC_OUT0[5]
    PORT
      LAYER met2 ;
        RECT 920.050 1044.980 1036.350 1045.760 ;
    END
  END ADC_OUT0[5]
  PIN ADC_OUT1[5]
    PORT
      LAYER met2 ;
        RECT 921.105 1062.070 1036.625 1062.980 ;
    END
  END ADC_OUT1[5]
  PIN ADC_OUT2[5]
    PORT
      LAYER met2 ;
        RECT 919.660 1080.690 1036.900 1081.450 ;
    END
  END ADC_OUT2[5]
  PIN ADC_OUT0[6]
    PORT
      LAYER met2 ;
        RECT 920.910 1105.840 1037.170 1106.580 ;
    END
  END ADC_OUT0[6]
  PIN ADC_OUT1[6]
    PORT
      LAYER met2 ;
        RECT 920.700 1122.810 1036.660 1123.610 ;
    END
  END ADC_OUT1[6]
  PIN ADC_OUT2[6]
    PORT
      LAYER met2 ;
        RECT 919.325 1141.420 1037.345 1142.250 ;
    END
  END ADC_OUT2[6]
  PIN ADC_OUT0[7]
    PORT
      LAYER met2 ;
        RECT 919.735 1166.560 1037.035 1167.410 ;
    END
  END ADC_OUT0[7]
  PIN ADC_OUT1[7]
    PORT
      LAYER met2 ;
        RECT 921.175 1183.640 1036.335 1184.450 ;
    END
  END ADC_OUT1[7]
  PIN ADC_OUT2[7]
    PORT
      LAYER met2 ;
        RECT 921.340 1202.160 1036.600 1203.040 ;
    END
  END ADC_OUT2[7]
  PIN ADC_OUT0[8]
    PORT
      LAYER met3 ;
        RECT 841.380 805.040 1036.070 806.000 ;
    END
  END ADC_OUT0[8]
  PIN ADC_OUT1[8]
    PORT
      LAYER met3 ;
        RECT 841.400 822.140 1036.420 823.100 ;
    END
  END ADC_OUT1[8]
  PIN ADC_OUT2[8]
    PORT
      LAYER met3 ;
        RECT 841.400 840.770 1036.800 841.730 ;
    END
  END ADC_OUT2[8]
  PIN ADC_OUT0[9]
    PORT
      LAYER met3 ;
        RECT 841.500 865.860 1036.340 866.820 ;
    END
  END ADC_OUT0[9]
  PIN ADC_OUT1[9]
    PORT
      LAYER met3 ;
        RECT 841.340 882.960 1036.000 883.920 ;
    END
  END ADC_OUT1[9]
  PIN ADC_OUT2[9]
    PORT
      LAYER met3 ;
        RECT 841.320 901.380 1036.310 902.340 ;
    END
  END ADC_OUT2[9]
  PIN ADC_OUT0[10]
    PORT
      LAYER met3 ;
        RECT 841.500 926.520 1036.210 927.480 ;
    END
  END ADC_OUT0[10]
  PIN ADC_OUT1[10]
    PORT
      LAYER met3 ;
        RECT 841.450 943.620 1036.000 944.580 ;
    END
  END ADC_OUT1[10]
  PIN ADC_OUT2[10]
    PORT
      LAYER met3 ;
        RECT 841.510 962.200 1035.560 963.160 ;
    END
  END ADC_OUT2[10]
  PIN ADC_OUT0[11]
    PORT
      LAYER met3 ;
        RECT 841.430 987.310 1036.640 988.270 ;
    END
  END ADC_OUT0[11]
  PIN ADC_OUT1[11]
    PORT
      LAYER met3 ;
        RECT 841.430 1004.350 1036.500 1005.310 ;
    END
  END ADC_OUT1[11]
  PIN ADC_OUT2[11]
    PORT
      LAYER met3 ;
        RECT 841.370 1023.020 1035.670 1023.980 ;
    END
  END ADC_OUT2[11]
  PIN ADC_OUT0[12]
    PORT
      LAYER met3 ;
        RECT 841.490 1048.190 1036.680 1049.150 ;
    END
  END ADC_OUT0[12]
  PIN ADC_OUT1[12]
    PORT
      LAYER met3 ;
        RECT 841.300 1065.110 1036.880 1066.070 ;
    END
  END ADC_OUT1[12]
  PIN ADC_OUT2[12]
    PORT
      LAYER met3 ;
        RECT 841.370 1083.690 1036.210 1084.650 ;
    END
  END ADC_OUT2[12]
  PIN ADC_OUT0[13]
    PORT
      LAYER met3 ;
        RECT 841.310 1108.740 1036.590 1109.700 ;
    END
  END ADC_OUT0[13]
  PIN ADC_OUT1[13]
    PORT
      LAYER met3 ;
        RECT 841.390 1125.930 1036.820 1126.890 ;
    END
  END ADC_OUT1[13]
  PIN ADC_OUT2[13]
    PORT
      LAYER met3 ;
        RECT 841.370 1144.410 1036.750 1145.370 ;
    END
  END ADC_OUT2[13]
  PIN ADC_OUT0[14]
    PORT
      LAYER met3 ;
        RECT 841.460 1169.620 1037.090 1170.580 ;
    END
  END ADC_OUT0[14]
  PIN ADC_OUT1[14]
    PORT
      LAYER met3 ;
        RECT 841.390 1186.630 1037.140 1187.590 ;
    END
  END ADC_OUT1[14]
  PIN ADC_OUT2[14]
    PORT
      LAYER met3 ;
        RECT 841.360 1205.170 1036.720 1206.130 ;
    END
  END ADC_OUT2[14]
  PIN ADC_OUT0[15]
    PORT
      LAYER met3 ;
        RECT 841.430 1230.380 1036.770 1231.340 ;
    END
  END ADC_OUT0[15]
  PIN ADC_OUT1[15]
    PORT
      LAYER met3 ;
        RECT 841.390 1247.430 1037.280 1248.390 ;
    END
  END ADC_OUT1[15]
  PIN ADC_OUT2[15]
    PORT
      LAYER met3 ;
        RECT 841.390 1266.050 1037.620 1267.010 ;
    END
  END ADC_OUT2[15]
  PIN PRE
    PORT
      LAYER met3 ;
        RECT 412.105 485.545 1033.695 486.515 ;
    END
  END PRE
  PIN CLK_EN_ADC[0]
    PORT
      LAYER met1 ;
        RECT 1022.865 1223.400 1039.390 1226.080 ;
    END
  END CLK_EN_ADC[0]
  PIN CLK_EN_ADC[1]
    PORT
      LAYER met1 ;
        RECT 1024.195 1283.770 1041.160 1286.370 ;
    END
  END CLK_EN_ADC[1]
  PIN REF_CSA
    PORT
      LAYER met2 ;
        RECT 612.745 730.000 615.475 1315.555 ;
    END
  END REF_CSA
  PIN SAEN_CSA
    PORT
      LAYER met1 ;
        RECT 856.395 509.840 1036.910 511.100 ;
    END
  END SAEN_CSA
  OBS
      LAYER li1 ;
        RECT -4.105 7.760 1033.835 1286.895 ;
      LAYER met1 ;
        RECT -3.650 1286.650 1033.830 1308.090 ;
        RECT -3.650 1283.490 1023.915 1286.650 ;
        RECT -3.650 1226.360 1033.830 1283.490 ;
        RECT -3.650 1223.120 1022.585 1226.360 ;
        RECT -3.650 511.380 1033.830 1223.120 ;
        RECT -3.650 509.560 856.115 511.380 ;
        RECT -3.650 8.215 1033.830 509.560 ;
      LAYER met2 ;
        RECT -10.490 729.720 612.465 1312.290 ;
        RECT 615.755 1312.015 1029.230 1312.290 ;
        RECT 615.755 1311.755 817.520 1312.015 ;
        RECT 615.755 1291.460 801.850 1311.755 ;
        RECT 803.920 1311.655 817.520 1311.755 ;
        RECT 803.920 1300.220 810.850 1311.655 ;
        RECT 813.080 1307.490 817.520 1311.655 ;
        RECT 819.650 1307.490 1029.230 1312.015 ;
        RECT 813.080 1300.220 1029.230 1307.490 ;
        RECT 803.920 1291.460 1029.230 1300.220 ;
        RECT 615.755 1203.320 1029.230 1291.460 ;
        RECT 615.755 1201.880 921.060 1203.320 ;
        RECT 615.755 1184.730 1029.230 1201.880 ;
        RECT 615.755 1183.360 920.895 1184.730 ;
        RECT 615.755 1167.690 1029.230 1183.360 ;
        RECT 615.755 1166.280 919.455 1167.690 ;
        RECT 615.755 1142.530 1029.230 1166.280 ;
        RECT 615.755 1141.140 919.045 1142.530 ;
        RECT 615.755 1123.890 1029.230 1141.140 ;
        RECT 615.755 1122.530 920.420 1123.890 ;
        RECT 615.755 1106.860 1029.230 1122.530 ;
        RECT 615.755 1105.560 920.630 1106.860 ;
        RECT 615.755 1081.730 1029.230 1105.560 ;
        RECT 615.755 1080.410 919.380 1081.730 ;
        RECT 615.755 1063.260 1029.230 1080.410 ;
        RECT 615.755 1061.790 920.825 1063.260 ;
        RECT 615.755 1046.040 1029.230 1061.790 ;
        RECT 615.755 1044.700 919.770 1046.040 ;
        RECT 615.755 1021.010 1029.230 1044.700 ;
        RECT 615.755 1019.650 919.690 1021.010 ;
        RECT 615.755 1002.430 1029.230 1019.650 ;
        RECT 615.755 1001.060 920.850 1002.430 ;
        RECT 615.755 985.400 1029.230 1001.060 ;
        RECT 615.755 984.030 920.745 985.400 ;
        RECT 615.755 960.310 1029.230 984.030 ;
        RECT 615.755 958.890 919.160 960.310 ;
        RECT 615.755 941.750 1029.230 958.890 ;
        RECT 615.755 940.290 920.130 941.750 ;
        RECT 615.755 924.660 1029.230 940.290 ;
        RECT 615.755 923.220 920.650 924.660 ;
        RECT 615.755 899.450 1029.230 923.220 ;
        RECT 615.755 898.080 919.565 899.450 ;
        RECT 615.755 880.880 1029.230 898.080 ;
        RECT 615.755 879.480 919.780 880.880 ;
        RECT 615.755 863.890 1029.230 879.480 ;
        RECT 615.755 862.470 919.510 863.890 ;
        RECT 615.755 838.750 1029.230 862.470 ;
        RECT 615.755 837.330 920.750 838.750 ;
        RECT 615.755 820.170 1029.230 837.330 ;
        RECT 615.755 818.750 920.730 820.170 ;
        RECT 615.755 803.050 1029.230 818.750 ;
        RECT 615.755 801.740 919.155 803.050 ;
        RECT 615.755 777.890 1029.230 801.740 ;
        RECT 615.755 776.570 919.550 777.890 ;
        RECT 615.755 759.350 1029.230 776.570 ;
        RECT 615.755 758.060 920.835 759.350 ;
        RECT 615.755 742.330 1029.230 758.060 ;
        RECT 615.755 740.960 920.890 742.330 ;
        RECT 615.755 729.720 1029.230 740.960 ;
        RECT -10.490 715.925 1029.230 729.720 ;
        RECT -10.490 714.475 750.715 715.925 ;
        RECT -10.490 702.905 1029.230 714.475 ;
        RECT -10.490 701.455 750.715 702.905 ;
        RECT -10.490 689.675 1029.230 701.455 ;
        RECT -10.490 688.225 750.715 689.675 ;
        RECT -10.490 676.565 1029.230 688.225 ;
        RECT -10.490 675.115 750.715 676.565 ;
        RECT -10.490 663.335 1029.230 675.115 ;
        RECT -10.490 661.885 750.715 663.335 ;
        RECT -10.490 650.265 1029.230 661.885 ;
        RECT -10.490 648.815 750.715 650.265 ;
        RECT -10.490 636.985 1029.230 648.815 ;
        RECT -10.490 635.535 750.715 636.985 ;
        RECT -10.490 623.905 1029.230 635.535 ;
        RECT -10.490 622.455 750.715 623.905 ;
        RECT -10.490 610.695 1029.230 622.455 ;
        RECT -10.490 609.245 750.715 610.695 ;
        RECT -10.490 597.605 1029.230 609.245 ;
        RECT -10.490 596.155 750.715 597.605 ;
        RECT -10.490 584.435 1029.230 596.155 ;
        RECT -10.490 582.985 750.715 584.435 ;
        RECT -10.490 571.225 1029.230 582.985 ;
        RECT -10.490 569.775 750.715 571.225 ;
        RECT -10.490 558.115 1029.230 569.775 ;
        RECT -10.490 556.665 750.715 558.115 ;
        RECT -10.490 544.965 1029.230 556.665 ;
        RECT -10.490 543.515 750.715 544.965 ;
        RECT -10.490 531.745 1029.230 543.515 ;
        RECT -10.490 530.295 750.715 531.745 ;
        RECT -10.490 518.595 1029.230 530.295 ;
        RECT -10.490 517.255 750.715 518.595 ;
        RECT -10.490 211.290 1029.230 517.255 ;
        RECT -10.490 211.070 437.780 211.290 ;
        RECT -10.490 -19.490 417.360 211.070 ;
        RECT 419.990 -19.490 437.780 211.070 ;
        RECT 440.610 211.270 1029.230 211.290 ;
        RECT 440.610 211.260 450.450 211.270 ;
        RECT 440.610 -19.490 441.210 211.260 ;
        RECT -10.490 -19.570 441.210 -19.490 ;
        RECT 444.040 -16.570 450.450 211.260 ;
        RECT 444.040 -19.570 445.230 -16.570 ;
        RECT 448.090 -19.490 450.450 -16.570 ;
        RECT 453.280 -19.490 1029.230 211.270 ;
        RECT 448.090 -19.570 1029.230 -19.490 ;
        RECT -10.490 -20.140 1029.230 -19.570 ;
      LAYER met3 ;
        RECT -30.190 927.045 -10.910 1315.590 ;
      LAYER met3 ;
        RECT -8.080 927.045 9.670 1315.590 ;
      LAYER met3 ;
        RECT -30.190 926.825 9.670 927.045 ;
      LAYER met3 ;
        RECT 12.270 1315.455 17.135 1315.590 ;
        RECT 12.270 926.855 13.025 1315.455 ;
        RECT 15.890 926.935 17.135 1315.455 ;
        RECT 20.000 1315.585 37.300 1315.590 ;
        RECT 20.000 926.935 22.225 1315.585 ;
        RECT 15.890 926.855 22.225 926.935 ;
        RECT 12.270 926.845 22.225 926.855 ;
        RECT 25.090 926.845 37.300 1315.585 ;
        RECT 12.270 926.825 37.300 926.845 ;
      LAYER met3 ;
        RECT -30.190 926.735 37.300 926.825 ;
      LAYER met3 ;
        RECT 40.700 926.785 50.370 1315.590 ;
        RECT 53.770 926.785 88.700 1315.590 ;
        RECT 40.700 926.775 88.700 926.785 ;
        RECT 92.100 1315.560 107.940 1315.590 ;
        RECT 92.100 926.795 101.860 1315.560 ;
        RECT 105.260 926.825 107.940 1315.560 ;
        RECT 111.340 926.865 121.020 1315.590 ;
        RECT 124.420 926.865 159.290 1315.590 ;
        RECT 111.340 926.825 159.290 926.865 ;
        RECT 105.260 926.795 159.290 926.825 ;
        RECT 92.100 926.785 159.290 926.795 ;
        RECT 162.690 1315.460 178.490 1315.590 ;
        RECT 162.690 926.835 172.380 1315.460 ;
        RECT 175.780 926.895 178.490 1315.460 ;
        RECT 181.890 926.895 191.570 1315.590 ;
        RECT 175.780 926.835 191.570 926.895 ;
        RECT 162.690 926.785 191.570 926.835 ;
        RECT 92.100 926.775 191.570 926.785 ;
        RECT 40.700 926.745 191.570 926.775 ;
        RECT 194.970 926.945 229.880 1315.590 ;
        RECT 233.280 1315.490 249.080 1315.590 ;
        RECT 233.280 926.945 243.030 1315.490 ;
        RECT 194.970 926.755 243.030 926.945 ;
        RECT 246.430 926.855 249.080 1315.490 ;
        RECT 252.480 926.895 262.130 1315.590 ;
        RECT 265.530 926.895 300.430 1315.590 ;
        RECT 252.480 926.855 300.430 926.895 ;
        RECT 303.830 926.855 313.450 1315.590 ;
        RECT 316.850 926.855 319.630 1315.590 ;
        RECT 246.430 926.815 319.630 926.855 ;
        RECT 323.030 1315.520 371.230 1315.590 ;
        RECT 323.030 926.815 332.790 1315.520 ;
        RECT 246.430 926.755 332.790 926.815 ;
        RECT 194.970 926.745 332.790 926.755 ;
        RECT 336.190 926.815 371.230 1315.520 ;
        RECT 374.630 926.855 384.370 1315.590 ;
        RECT 387.770 926.855 390.430 1315.590 ;
        RECT 374.630 926.815 390.430 926.855 ;
        RECT 393.830 926.895 403.500 1315.590 ;
        RECT 406.900 926.895 441.850 1315.590 ;
        RECT 393.830 926.815 441.850 926.895 ;
        RECT 336.190 926.775 441.850 926.815 ;
        RECT 445.250 927.025 454.970 1315.590 ;
        RECT 458.370 927.025 460.890 1315.590 ;
        RECT 445.250 926.945 460.890 927.025 ;
        RECT 464.290 926.945 473.970 1315.590 ;
        RECT 445.250 926.815 473.970 926.945 ;
        RECT 477.370 926.945 512.470 1315.590 ;
        RECT 515.870 926.945 525.270 1315.590 ;
        RECT 477.370 926.895 525.270 926.945 ;
        RECT 528.670 926.895 531.560 1315.590 ;
        RECT 477.370 926.815 531.560 926.895 ;
        RECT 534.960 926.945 544.590 1315.590 ;
        RECT 547.990 926.945 582.990 1315.590 ;
        RECT 534.960 926.895 582.990 926.945 ;
        RECT 586.390 1311.990 596.160 1315.590 ;
        RECT 599.870 1311.990 1029.205 1315.590 ;
        RECT 586.390 1267.410 1029.205 1311.990 ;
        RECT 586.390 1265.650 840.990 1267.410 ;
        RECT 586.390 1248.790 1029.205 1265.650 ;
        RECT 586.390 1247.030 840.990 1248.790 ;
        RECT 586.390 1231.740 1029.205 1247.030 ;
        RECT 586.390 1229.980 841.030 1231.740 ;
        RECT 586.390 1206.530 1029.205 1229.980 ;
        RECT 586.390 1204.770 840.960 1206.530 ;
        RECT 586.390 1187.990 1029.205 1204.770 ;
        RECT 586.390 1186.230 840.990 1187.990 ;
        RECT 586.390 1170.980 1029.205 1186.230 ;
        RECT 586.390 1169.220 841.060 1170.980 ;
        RECT 586.390 1145.770 1029.205 1169.220 ;
        RECT 586.390 1144.010 840.970 1145.770 ;
        RECT 586.390 1127.290 1029.205 1144.010 ;
        RECT 586.390 1125.530 840.990 1127.290 ;
        RECT 586.390 1110.100 1029.205 1125.530 ;
        RECT 586.390 1108.340 840.910 1110.100 ;
        RECT 586.390 1085.050 1029.205 1108.340 ;
        RECT 586.390 1083.290 840.970 1085.050 ;
        RECT 586.390 1066.470 1029.205 1083.290 ;
        RECT 586.390 1064.710 840.900 1066.470 ;
        RECT 586.390 1049.550 1029.205 1064.710 ;
        RECT 586.390 1047.790 841.090 1049.550 ;
        RECT 586.390 1024.380 1029.205 1047.790 ;
        RECT 586.390 1022.620 840.970 1024.380 ;
        RECT 586.390 1005.710 1029.205 1022.620 ;
        RECT 586.390 1003.950 841.030 1005.710 ;
        RECT 586.390 988.670 1029.205 1003.950 ;
        RECT 586.390 986.910 841.030 988.670 ;
        RECT 586.390 963.560 1029.205 986.910 ;
        RECT 586.390 961.800 841.110 963.560 ;
        RECT 586.390 944.980 1029.205 961.800 ;
        RECT 586.390 943.220 841.050 944.980 ;
        RECT 586.390 927.880 1029.205 943.220 ;
        RECT 586.390 926.895 841.100 927.880 ;
        RECT 534.960 926.815 841.100 926.895 ;
        RECT 445.250 926.775 841.100 926.815 ;
        RECT 336.190 926.745 841.100 926.775 ;
        RECT 40.700 926.735 841.100 926.745 ;
      LAYER met3 ;
        RECT -30.190 926.120 841.100 926.735 ;
        RECT -30.190 902.740 1029.205 926.120 ;
        RECT -30.190 900.980 840.920 902.740 ;
        RECT -30.190 884.320 1029.205 900.980 ;
        RECT -30.190 882.560 840.940 884.320 ;
        RECT -30.190 867.220 1029.205 882.560 ;
        RECT -30.190 865.460 841.100 867.220 ;
        RECT -30.190 842.130 1029.205 865.460 ;
        RECT -30.190 840.370 841.000 842.130 ;
        RECT -30.190 823.500 1029.205 840.370 ;
        RECT -30.190 821.740 841.000 823.500 ;
        RECT -30.190 806.400 1029.205 821.740 ;
        RECT -30.190 804.640 840.980 806.400 ;
        RECT -30.190 729.540 1029.205 804.640 ;
        RECT -30.190 725.040 782.655 729.540 ;
        RECT -30.190 611.530 1029.205 725.040 ;
      LAYER met3 ;
        RECT 0.535 608.080 1029.205 611.530 ;
      LAYER met3 ;
        RECT -30.190 598.320 1029.205 608.080 ;
      LAYER met3 ;
        RECT 0.495 594.870 1029.205 598.320 ;
      LAYER met3 ;
        RECT -30.190 559.920 1029.205 594.870 ;
      LAYER met3 ;
        RECT 0.445 556.470 1029.205 559.920 ;
      LAYER met3 ;
        RECT -30.190 546.840 1029.205 556.470 ;
      LAYER met3 ;
        RECT 0.575 543.390 1029.205 546.840 ;
      LAYER met3 ;
        RECT -30.190 540.650 1029.205 543.390 ;
      LAYER met3 ;
        RECT 0.495 537.200 1029.205 540.650 ;
      LAYER met3 ;
        RECT -30.190 527.750 1029.205 537.200 ;
      LAYER met3 ;
        RECT -26.880 524.250 1029.205 527.750 ;
      LAYER met3 ;
        RECT -30.190 489.240 1029.205 524.250 ;
      LAYER met3 ;
        RECT 0.575 486.915 1029.205 489.240 ;
        RECT 0.575 485.790 411.705 486.915 ;
      LAYER met3 ;
        RECT -30.190 485.145 411.705 485.790 ;
        RECT -30.190 476.190 1029.205 485.145 ;
      LAYER met3 ;
        RECT 0.445 472.740 1029.205 476.190 ;
      LAYER met3 ;
        RECT -30.190 470.100 1029.205 472.740 ;
      LAYER met3 ;
        RECT 0.365 466.650 1029.205 470.100 ;
      LAYER met3 ;
        RECT -30.190 457.070 1029.205 466.650 ;
      LAYER met3 ;
        RECT 0.615 453.620 1029.205 457.070 ;
      LAYER met3 ;
        RECT -30.190 418.590 1029.205 453.620 ;
      LAYER met3 ;
        RECT 0.495 415.140 1029.205 418.590 ;
      LAYER met3 ;
        RECT -30.190 405.710 1029.205 415.140 ;
      LAYER met3 ;
        RECT 0.575 402.260 1029.205 405.710 ;
      LAYER met3 ;
        RECT -30.190 399.480 1029.205 402.260 ;
      LAYER met3 ;
        RECT 0.535 396.030 1029.205 399.480 ;
      LAYER met3 ;
        RECT -30.190 386.470 1029.205 396.030 ;
      LAYER met3 ;
        RECT 0.575 383.020 1029.205 386.470 ;
      LAYER met3 ;
        RECT -30.190 348.120 1029.205 383.020 ;
      LAYER met3 ;
        RECT 0.645 344.670 1029.205 348.120 ;
      LAYER met3 ;
        RECT -30.190 334.860 1029.205 344.670 ;
      LAYER met3 ;
        RECT 0.575 331.410 1029.205 334.860 ;
      LAYER met3 ;
        RECT -30.190 328.780 1029.205 331.410 ;
      LAYER met3 ;
        RECT 0.535 325.330 1029.205 328.780 ;
      LAYER met3 ;
        RECT -30.190 315.870 1029.205 325.330 ;
      LAYER met3 ;
        RECT -26.830 312.370 1029.205 315.870 ;
      LAYER met3 ;
        RECT -30.190 277.440 1029.205 312.370 ;
      LAYER met3 ;
        RECT 0.495 273.990 1029.205 277.440 ;
      LAYER met3 ;
        RECT -30.190 264.260 1029.205 273.990 ;
      LAYER met3 ;
        RECT 0.535 260.810 1029.205 264.260 ;
      LAYER met3 ;
        RECT -30.190 258.200 1029.205 260.810 ;
        RECT -30.190 254.700 -30.140 258.200 ;
      LAYER met3 ;
        RECT -26.690 254.700 1029.205 258.200 ;
      LAYER met3 ;
        RECT -30.190 245.150 1029.205 254.700 ;
      LAYER met3 ;
        RECT 0.445 241.700 1029.205 245.150 ;
      LAYER met3 ;
        RECT -30.190 211.500 1029.205 241.700 ;
        RECT -30.190 206.640 465.530 211.500 ;
        RECT -30.190 203.190 -30.140 206.640 ;
      LAYER met3 ;
        RECT 0.645 203.190 465.530 206.640 ;
      LAYER met3 ;
        RECT -30.190 193.730 465.530 203.190 ;
      LAYER met3 ;
        RECT 0.495 190.280 465.530 193.730 ;
      LAYER met3 ;
        RECT -30.190 187.730 465.530 190.280 ;
      LAYER met3 ;
        RECT 0.555 184.280 465.530 187.730 ;
      LAYER met3 ;
        RECT -30.190 174.550 465.530 184.280 ;
      LAYER met3 ;
        RECT 0.605 171.100 465.530 174.550 ;
      LAYER met3 ;
        RECT -30.190 136.310 465.530 171.100 ;
      LAYER met3 ;
        RECT 0.525 132.860 465.530 136.310 ;
      LAYER met3 ;
        RECT -30.190 123.210 465.530 132.860 ;
        RECT -30.190 119.760 -30.160 123.210 ;
      LAYER met3 ;
        RECT 0.565 119.760 465.530 123.210 ;
      LAYER met3 ;
        RECT -30.190 117.150 465.530 119.760 ;
        RECT -30.190 113.650 -30.160 117.150 ;
      LAYER met3 ;
        RECT -26.710 113.650 465.530 117.150 ;
      LAYER met3 ;
        RECT -30.190 104.020 465.530 113.650 ;
      LAYER met3 ;
        RECT 0.615 100.570 465.530 104.020 ;
      LAYER met3 ;
        RECT -30.190 65.610 465.530 100.570 ;
        RECT -30.190 62.160 -30.180 65.610 ;
      LAYER met3 ;
        RECT 0.605 62.160 465.530 65.610 ;
      LAYER met3 ;
        RECT -30.190 52.570 465.530 62.160 ;
        RECT -30.190 49.120 -30.150 52.570 ;
      LAYER met3 ;
        RECT 0.655 49.120 465.530 52.570 ;
      LAYER met3 ;
        RECT -30.190 36.930 465.530 49.120 ;
      LAYER met3 ;
        RECT 0.545 33.910 465.530 36.930 ;
      LAYER met3 ;
        RECT -30.190 31.730 465.530 33.910 ;
      LAYER met3 ;
        RECT 0.455 28.900 465.530 31.730 ;
      LAYER met3 ;
        RECT -30.190 27.560 465.530 28.900 ;
      LAYER met3 ;
        RECT 0.535 24.730 465.530 27.560 ;
      LAYER met3 ;
        RECT -30.190 24.210 465.530 24.730 ;
      LAYER met3 ;
        RECT 0.565 21.380 465.530 24.210 ;
      LAYER met3 ;
        RECT -30.190 3.775 465.530 21.380 ;
      LAYER met3 ;
        RECT 0.345 0.945 465.530 3.775 ;
      LAYER met3 ;
        RECT -30.190 -19.170 465.530 0.945 ;
      LAYER met3 ;
        RECT 469.100 211.490 1029.205 211.500 ;
        RECT 469.100 211.460 619.740 211.490 ;
        RECT 469.100 211.450 516.790 211.460 ;
        RECT 469.100 -19.170 478.570 211.450 ;
        RECT 482.140 -19.170 516.790 211.450 ;
        RECT 520.360 211.450 619.740 211.460 ;
        RECT 520.360 211.440 587.400 211.450 ;
        RECT 520.360 -19.170 529.920 211.440 ;
        RECT 533.490 211.410 587.400 211.440 ;
        RECT 533.490 -19.170 536.170 211.410 ;
        RECT 539.740 211.370 587.400 211.410 ;
        RECT 539.740 -19.170 549.260 211.370 ;
        RECT 552.830 -19.170 587.400 211.370 ;
        RECT 590.970 211.400 619.740 211.450 ;
        RECT 590.970 -19.170 600.560 211.400 ;
        RECT 604.130 211.340 619.740 211.400 ;
        RECT 604.130 -19.170 606.360 211.340 ;
        RECT 609.930 -19.170 619.740 211.340 ;
        RECT 623.310 211.480 760.860 211.490 ;
        RECT 623.310 211.290 670.960 211.480 ;
        RECT 623.310 -19.170 657.960 211.290 ;
        RECT 661.530 -19.170 670.960 211.290 ;
        RECT 674.530 211.420 760.860 211.480 ;
        RECT 674.530 211.380 747.700 211.420 ;
        RECT 674.530 211.340 728.560 211.380 ;
        RECT 674.530 170.345 690.300 211.340 ;
        RECT 674.530 -19.170 677.210 170.345 ;
        RECT 680.780 -19.170 690.300 170.345 ;
        RECT 693.870 -19.170 728.560 211.340 ;
        RECT 732.130 -19.170 741.400 211.380 ;
        RECT 744.970 -19.170 747.700 211.380 ;
        RECT 751.270 -19.170 760.860 211.420 ;
        RECT 764.430 211.460 1029.205 211.490 ;
        RECT 764.430 211.420 869.980 211.460 ;
        RECT 764.430 -19.170 799.380 211.420 ;
        RECT 802.950 211.380 818.420 211.420 ;
        RECT 802.950 -19.170 812.420 211.380 ;
        RECT 815.990 -19.170 818.420 211.380 ;
        RECT 821.990 211.340 869.980 211.420 ;
        RECT 821.990 -19.160 831.550 211.340 ;
        RECT 835.120 -19.160 869.980 211.340 ;
        RECT 821.990 -19.170 869.980 -19.160 ;
        RECT 873.550 211.420 1029.205 211.460 ;
        RECT 873.550 211.290 902.160 211.420 ;
        RECT 873.550 211.210 889.070 211.290 ;
        RECT 873.550 -19.170 882.980 211.210 ;
        RECT 886.550 -19.170 889.070 211.210 ;
        RECT 892.640 -19.170 902.160 211.290 ;
        RECT 905.730 211.340 959.670 211.420 ;
        RECT 905.730 211.290 953.705 211.340 ;
        RECT 905.730 -19.170 940.540 211.290 ;
        RECT 944.110 -19.170 953.705 211.290 ;
        RECT 957.115 -19.170 959.670 211.340 ;
        RECT 963.240 211.380 1029.205 211.420 ;
        RECT 963.240 211.340 1024.400 211.380 ;
        RECT 963.240 211.290 1011.270 211.340 ;
        RECT 963.240 -19.170 972.720 211.290 ;
        RECT 976.290 -19.170 1011.270 211.290 ;
        RECT 1014.840 -19.170 1024.400 211.340 ;
        RECT 1027.970 -19.170 1029.205 211.380 ;
  END
END RRAM_ANALOG
END LIBRARY

